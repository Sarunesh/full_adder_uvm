`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "fa_common.sv"
`include "fa_interface.sv"
`include "full_adder.v"
`include "fa_tx.sv"
`include "fa_seq_lib.sv"
`include "fa_sqr.sv"
`include "fa_drv.sv"
`include "fa_mon.sv"
`include "fa_sub.sv"
`include "fa_sbd.sv"
`include "fa_agent.sv"
`include "fa_env.sv"
`include "test_lib.sv"
`include "top.sv"
