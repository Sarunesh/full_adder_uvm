typedef uvm_sequencer#(fa_tx) fa_sqr;
