interface fa_interface(input reg rst);
	logic sum;
	logic carry;
	logic a;
	logic b;
	logic cin;	
endinterface
